module apb_slave(apb_interface apb_if);

    // Device registers
    logic [31:0] data_reg;      // Data register (value to add)
    logic [1:0] control_reg;   // Control register
    logic [31:0] result_reg;    // Result register (current accumulated result)

    // Register address definitions
    localparam DATA_ADDR    = 8'h00;  
    localparam CONTROL_ADDR = 8'h04;   
    localparam RESULT_ADDR  = 8'h08;  

    // Control register bits
    localparam START_BIT = 0;  // bit 0 - start OR accumulation
    localparam RESET_BIT = 1;  // bit 1 - reset result register

    always_ff @(posedge apb_if.PCLK or negedge apb_if.PRESETn) begin
        if (!apb_if.PRESETn) begin
            // Reset registers
            data_reg <= 32'h0;
            control_reg <= 2'b00;    
            result_reg <= 32'h0;
            apb_if.PREADY <= 1'b0;
            apb_if.PSLVERR <= 1'b0;
            apb_if.PRDATA <= 32'h0;
        end
        else begin
            apb_if.PSLVERR <= 1'b0;
            apb_if.PREADY <= 1'b0;
            
            // Write operations
            if (apb_if.PSEL && apb_if.PENABLE && apb_if.PWRITE) begin
                apb_if.PREADY <= 1'b1;
                
                case (apb_if.PADDR)
                    DATA_ADDR: begin
                        data_reg <= apb_if.PWDATA;
                        if(!apb_if.PREADY) $display("[APB_SLAVE] Write DATA register: %h", apb_if.PWDATA);
                    end
                    CONTROL_ADDR: begin
                        control_reg <= apb_if.PWDATA[1:0]; 
                        if(!apb_if.PREADY) $display("[APB_SLAVE] Write CONTROL register: %b", apb_if.PWDATA[1:0]);
                        
                        // Reset result register if reset bit is set
                        if (apb_if.PWDATA[RESET_BIT]) begin
                            result_reg <= 32'h0;
                            if(!apb_if.PREADY) $display("[APB_SLAVE] Reset result register");
                        end
                        // OR accumulation if start bit is set (and not resetting)
                        else if (apb_if.PWDATA[START_BIT]) begin
                            result_reg <= result_reg | data_reg;
                            if(!apb_if.PREADY) $display("[APB_SLAVE] OR accumulation: result = %h", result_reg | data_reg);
                        end
                    end
                    RESULT_ADDR: begin
                        // Result register is read-only - error on write attempt
                        apb_if.PSLVERR <= 1'b1;
                        if(!apb_if.PREADY) $display("[APB_SLAVE] ERROR: Attempt to write to read-only RESULT register");
                    end
                    default: begin
                        apb_if.PSLVERR <= 1'b1;
                        if(!apb_if.PREADY) $display("[APB_SLAVE] ERROR: Invalid address %h", apb_if.PADDR);
                    end
                endcase
            end
            
            // Read operations
            else if (apb_if.PSEL && apb_if.PENABLE && !apb_if.PWRITE) begin
                apb_if.PREADY <= 1'b1;
                
                case (apb_if.PADDR)
                    DATA_ADDR: begin
                        apb_if.PRDATA <= data_reg;
                        if(!apb_if.PREADY) $display("[APB_SLAVE] Read DATA register: %h", data_reg);
                    end
                    CONTROL_ADDR: begin
                        apb_if.PRDATA <= {30'b0, control_reg}; 
                        if(!apb_if.PREADY) $display("[APB_SLAVE] Read CONTROL register: %b", control_reg);
                    end
                    RESULT_ADDR: begin
                        apb_if.PRDATA <= result_reg;
                        if(!apb_if.PREADY) $display("[APB_SLAVE] Read RESULT register: %h", result_reg);
                    end
                    default: begin
                        apb_if.PRDATA <= 32'h0;
                        apb_if.PSLVERR <= 1'b1;
                        if(!apb_if.PREADY) $display("[APB_SLAVE] ERROR: Invalid address %h", apb_if.PADDR);
                    end
                endcase
            end
        end
    end

endmodule
